
module soc_system (
	clk_clk,
	reset_reset_n,
	leds_0_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	leds_0_external_connection_export;
endmodule
