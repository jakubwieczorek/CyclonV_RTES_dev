// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		input  wire       clk_clk,                           //                        clk.clk
		output wire [7:0] leds_0_external_connection_export, // leds_0_external_connection.export
		input  wire       reset_reset_n                      //                      reset.reset_n
	);

	wire  [31:0] cpu_0_data_master_readdata;                                      // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_waitrequest;                                   // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire         cpu_0_data_master_debugaccess;                                   // cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire  [17:0] cpu_0_data_master_address;                                       // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;                                    // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_0_data_master_read;                                          // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire         cpu_0_data_master_readdatavalid;                                 // mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	wire         cpu_0_data_master_write;                                         // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                                     // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [31:0] cpu_1_data_master_readdata;                                      // mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_waitrequest;                                   // mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	wire         cpu_1_data_master_debugaccess;                                   // cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	wire  [17:0] cpu_1_data_master_address;                                       // cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	wire   [3:0] cpu_1_data_master_byteenable;                                    // cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	wire         cpu_1_data_master_read;                                          // cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	wire         cpu_1_data_master_readdatavalid;                                 // mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	wire         cpu_1_data_master_write;                                         // cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	wire  [31:0] cpu_1_data_master_writedata;                                     // cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	wire  [31:0] cpu_1_instruction_master_readdata;                               // mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	wire         cpu_1_instruction_master_waitrequest;                            // mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	wire  [17:0] cpu_1_instruction_master_address;                                // cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	wire         cpu_1_instruction_master_read;                                   // cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	wire         cpu_1_instruction_master_readdatavalid;                          // mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	wire  [31:0] cpu_0_instruction_master_readdata;                               // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;                            // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [17:0] cpu_0_instruction_master_address;                                // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                                   // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire         cpu_0_instruction_master_readdatavalid;                          // mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;        // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;     // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_interrupt_counter_0_avalon_slave_0_chipselect; // mm_interconnect_0:interrupt_counter_0_avalon_slave_0_chipselect -> interrupt_counter_0:ChipSelect
	wire  [31:0] mm_interconnect_0_interrupt_counter_0_avalon_slave_0_readdata;   // interrupt_counter_0:ReadData -> mm_interconnect_0:interrupt_counter_0_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_0_interrupt_counter_0_avalon_slave_0_address;    // mm_interconnect_0:interrupt_counter_0_avalon_slave_0_address -> interrupt_counter_0:Address
	wire         mm_interconnect_0_interrupt_counter_0_avalon_slave_0_read;       // mm_interconnect_0:interrupt_counter_0_avalon_slave_0_read -> interrupt_counter_0:Read
	wire         mm_interconnect_0_interrupt_counter_0_avalon_slave_0_write;      // mm_interconnect_0:interrupt_counter_0_avalon_slave_0_write -> interrupt_counter_0:Write
	wire  [31:0] mm_interconnect_0_interrupt_counter_0_avalon_slave_0_writedata;  // mm_interconnect_0:interrupt_counter_0_avalon_slave_0_writedata -> interrupt_counter_0:WriteData
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata;     // mailbox_simple_0:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_readdata
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest;  // mailbox_simple_0:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_waitrequest
	wire   [1:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address;      // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_address -> mailbox_simple_0:avmm_snd_address
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read;         // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_read -> mailbox_simple_0:avmm_snd_read
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write;        // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_write -> mailbox_simple_0:avmm_snd_write
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata;    // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_writedata -> mailbox_simple_0:avmm_snd_writedata
	wire  [31:0] mm_interconnect_0_perf_count_0_control_slave_readdata;           // perf_count_0:readdata -> mm_interconnect_0:perf_count_0_control_slave_readdata
	wire   [3:0] mm_interconnect_0_perf_count_0_control_slave_address;            // mm_interconnect_0:perf_count_0_control_slave_address -> perf_count_0:address
	wire         mm_interconnect_0_perf_count_0_control_slave_begintransfer;      // mm_interconnect_0:perf_count_0_control_slave_begintransfer -> perf_count_0:begintransfer
	wire         mm_interconnect_0_perf_count_0_control_slave_write;              // mm_interconnect_0:perf_count_0_control_slave_write -> perf_count_0:write
	wire  [31:0] mm_interconnect_0_perf_count_0_control_slave_writedata;          // mm_interconnect_0:perf_count_0_control_slave_writedata -> perf_count_0:writedata
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_readdata;                // cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest;             // cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess;             // mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_0_debug_mem_slave_address;                 // mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_read;                    // mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_0_debug_mem_slave_byteenable;              // mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_write;                   // mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_writedata;               // mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                  // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;                   // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                     // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                 // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                     // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_mutex_0_s1_chipselect;                         // mm_interconnect_0:mutex_0_s1_chipselect -> mutex_0:chipselect
	wire  [31:0] mm_interconnect_0_mutex_0_s1_readdata;                           // mutex_0:data_to_cpu -> mm_interconnect_0:mutex_0_s1_readdata
	wire   [0:0] mm_interconnect_0_mutex_0_s1_address;                            // mm_interconnect_0:mutex_0_s1_address -> mutex_0:address
	wire         mm_interconnect_0_mutex_0_s1_read;                               // mm_interconnect_0:mutex_0_s1_read -> mutex_0:read
	wire         mm_interconnect_0_mutex_0_s1_write;                              // mm_interconnect_0:mutex_0_s1_write -> mutex_0:write
	wire  [31:0] mm_interconnect_0_mutex_0_s1_writedata;                          // mm_interconnect_0:mutex_0_s1_writedata -> mutex_0:data_from_cpu
	wire         mm_interconnect_0_leds_0_s1_chipselect;                          // mm_interconnect_0:leds_0_s1_chipselect -> leds_0:chipselect
	wire  [31:0] mm_interconnect_0_leds_0_s1_readdata;                            // leds_0:readdata -> mm_interconnect_0:leds_0_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_0_s1_address;                             // mm_interconnect_0:leds_0_s1_address -> leds_0:address
	wire         mm_interconnect_0_leds_0_s1_write;                               // mm_interconnect_0:leds_0_s1_write -> leds_0:write_n
	wire  [31:0] mm_interconnect_0_leds_0_s1_writedata;                           // mm_interconnect_0:leds_0_s1_writedata -> leds_0:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                         // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                           // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                            // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                              // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                          // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata;        // jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest;     // jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> jtag_uart_1:av_read_n
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> jtag_uart_1:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata;   // mailbox_simple_0:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_readdata
	wire   [1:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address;    // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_address -> mailbox_simple_0:avmm_rcv_address
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read;       // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_read -> mailbox_simple_0:avmm_rcv_read
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write;      // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_write -> mailbox_simple_0:avmm_rcv_write
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata;  // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_writedata -> mailbox_simple_0:avmm_rcv_writedata
	wire  [31:0] mm_interconnect_0_perf_count_1_control_slave_readdata;           // perf_count_1:readdata -> mm_interconnect_0:perf_count_1_control_slave_readdata
	wire   [3:0] mm_interconnect_0_perf_count_1_control_slave_address;            // mm_interconnect_0:perf_count_1_control_slave_address -> perf_count_1:address
	wire         mm_interconnect_0_perf_count_1_control_slave_begintransfer;      // mm_interconnect_0:perf_count_1_control_slave_begintransfer -> perf_count_1:begintransfer
	wire         mm_interconnect_0_perf_count_1_control_slave_write;              // mm_interconnect_0:perf_count_1_control_slave_write -> perf_count_1:write
	wire  [31:0] mm_interconnect_0_perf_count_1_control_slave_writedata;          // mm_interconnect_0:perf_count_1_control_slave_writedata -> perf_count_1:writedata
	wire  [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_readdata;                // cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest;             // cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess;             // mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_1_debug_mem_slave_address;                 // mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_read;                    // mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_1_debug_mem_slave_byteenable;              // mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_write;                   // mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_writedata;               // mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;                // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;                  // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_1_s1_address;                   // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;                // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                     // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;                 // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                     // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire         mm_interconnect_0_timer_1_s1_chipselect;                         // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                           // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                            // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                              // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                          // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver2_irq;                                        // jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                        // timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_0_irq_irq;                                                   // irq_mapper:sender_irq -> cpu_0:irq
	wire         irq_mapper_001_receiver2_irq;                                    // jtag_uart_1:av_irq -> irq_mapper_001:receiver2_irq
	wire         irq_mapper_001_receiver3_irq;                                    // timer_1:irq -> irq_mapper_001:receiver3_irq
	wire  [31:0] cpu_1_irq_irq;                                                   // irq_mapper_001:sender_irq -> cpu_1:irq
	wire         irq_mapper_receiver1_irq;                                        // interrupt_counter_0:IRQ -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	wire         irq_mapper_receiver0_irq;                                        // mailbox_simple_0:irq_msg -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [cpu_0:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, perf_count_0:reset_n, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [cpu_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_0_debug_reset_request_reset;                                 // cpu_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in2]
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [cpu_1:reset_n, irq_mapper_001:reset, jtag_uart_1:rst_n, mm_interconnect_0:cpu_1_reset_reset_bridge_in_reset_reset, onchip_memory2_1:reset, perf_count_1:reset_n, rst_translator_001:in_reset, timer_1:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                          // rst_controller_001:reset_req -> [cpu_1:reset_req, onchip_memory2_1:reset_req, rst_translator_001:reset_req_in]
	wire         cpu_1_debug_reset_request_reset;                                 // cpu_1:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [interrupt_counter_0:nReset, leds_0:reset_n, mailbox_simple_0:rst_n, mm_interconnect_0:interrupt_counter_0_reset_sink_reset_bridge_in_reset_reset, mutex_0:reset_n]

	soc_system_cpu_0 cpu_0 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (cpu_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	soc_system_cpu_1 cpu_1 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (cpu_1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_1_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_1_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	counter interrupt_counter_0 (
		.Clk        (clk_clk),                                                         //            clock.clk
		.IRQ        (irq_mapper_receiver1_irq),                                        // interrupt_sender.irq
		.nReset     (~rst_controller_002_reset_out_reset),                             //       reset_sink.reset_n
		.Address    (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_address),    //   avalon_slave_0.address
		.ChipSelect (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_chipselect), //                 .chipselect
		.Read       (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_read),       //                 .read
		.Write      (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_write),      //                 .write
		.ReadData   (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_readdata),   //                 .readdata
		.WriteData  (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_writedata)   //                 .writedata
	);

	soc_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	soc_system_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver2_irq)                                 //               irq.irq
	);

	soc_system_leds_0 leds_0 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_leds_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_0_s1_readdata),   //                    .readdata
		.out_port   (leds_0_external_connection_export)       // external_connection.export
	);

	altera_avalon_mailbox #(
		.DWIDTH (32),
		.AWIDTH (2)
	) mailbox_simple_0 (
		.clk                  (clk_clk),                                                        //                   clk.clk
		.rst_n                (~rst_controller_002_reset_out_reset),                            //                 rst_n.reset_n
		.avmm_snd_address     (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address),     //       avmm_msg_sender.address
		.avmm_snd_writedata   (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata),   //                      .writedata
		.avmm_snd_write       (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write),       //                      .write
		.avmm_snd_read        (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read),        //                      .read
		.avmm_snd_readdata    (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata),    //                      .readdata
		.avmm_snd_waitrequest (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest), //                      .waitrequest
		.irq_msg              (irq_mapper_receiver0_irq),                                       // interrupt_msg_pending.irq
		.avmm_rcv_address     (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address),   //     avmm_msg_receiver.address
		.avmm_rcv_read        (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read),      //                      .read
		.avmm_rcv_writedata   (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata), //                      .writedata
		.avmm_rcv_write       (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write),     //                      .write
		.avmm_rcv_readdata    (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata),  //                      .readdata
		.irq_space            ()                                                                //           (terminated)
	);

	soc_system_mutex_0 mutex_0 (
		.reset_n       (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.clk           (clk_clk),                                 //   clk.clk
		.chipselect    (mm_interconnect_0_mutex_0_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_0_mutex_0_s1_writedata),  //      .writedata
		.read          (mm_interconnect_0_mutex_0_s1_read),       //      .read
		.write         (mm_interconnect_0_mutex_0_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_0_mutex_0_s1_readdata),   //      .readdata
		.address       (mm_interconnect_0_mutex_0_s1_address)     //      .address
	);

	soc_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_system_onchip_memory2_1 onchip_memory2_1 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_system_perf_count_0 perf_count_0 (
		.clk           (clk_clk),                                                    //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                            //         reset.reset_n
		.address       (mm_interconnect_0_perf_count_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_perf_count_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_perf_count_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_perf_count_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_perf_count_0_control_slave_writedata)      //              .writedata
	);

	soc_system_perf_count_0 perf_count_1 (
		.clk           (clk_clk),                                                    //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                        //         reset.reset_n
		.address       (mm_interconnect_0_perf_count_1_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_perf_count_1_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_perf_count_1_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_perf_count_1_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_perf_count_1_control_slave_writedata)      //              .writedata
	);

	soc_system_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	soc_system_timer_0 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver3_irq)             //   irq.irq
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                              (clk_clk),                                                         //                                            clk_0_clk.clk
		.cpu_0_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                                  //                    cpu_0_reset_reset_bridge_in_reset.reset
		.cpu_1_reset_reset_bridge_in_reset_reset                    (rst_controller_001_reset_out_reset),                              //                    cpu_1_reset_reset_bridge_in_reset.reset
		.interrupt_counter_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                              // interrupt_counter_0_reset_sink_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                                  (cpu_0_data_master_address),                                       //                                    cpu_0_data_master.address
		.cpu_0_data_master_waitrequest                              (cpu_0_data_master_waitrequest),                                   //                                                     .waitrequest
		.cpu_0_data_master_byteenable                               (cpu_0_data_master_byteenable),                                    //                                                     .byteenable
		.cpu_0_data_master_read                                     (cpu_0_data_master_read),                                          //                                                     .read
		.cpu_0_data_master_readdata                                 (cpu_0_data_master_readdata),                                      //                                                     .readdata
		.cpu_0_data_master_readdatavalid                            (cpu_0_data_master_readdatavalid),                                 //                                                     .readdatavalid
		.cpu_0_data_master_write                                    (cpu_0_data_master_write),                                         //                                                     .write
		.cpu_0_data_master_writedata                                (cpu_0_data_master_writedata),                                     //                                                     .writedata
		.cpu_0_data_master_debugaccess                              (cpu_0_data_master_debugaccess),                                   //                                                     .debugaccess
		.cpu_0_instruction_master_address                           (cpu_0_instruction_master_address),                                //                             cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest                       (cpu_0_instruction_master_waitrequest),                            //                                                     .waitrequest
		.cpu_0_instruction_master_read                              (cpu_0_instruction_master_read),                                   //                                                     .read
		.cpu_0_instruction_master_readdata                          (cpu_0_instruction_master_readdata),                               //                                                     .readdata
		.cpu_0_instruction_master_readdatavalid                     (cpu_0_instruction_master_readdatavalid),                          //                                                     .readdatavalid
		.cpu_1_data_master_address                                  (cpu_1_data_master_address),                                       //                                    cpu_1_data_master.address
		.cpu_1_data_master_waitrequest                              (cpu_1_data_master_waitrequest),                                   //                                                     .waitrequest
		.cpu_1_data_master_byteenable                               (cpu_1_data_master_byteenable),                                    //                                                     .byteenable
		.cpu_1_data_master_read                                     (cpu_1_data_master_read),                                          //                                                     .read
		.cpu_1_data_master_readdata                                 (cpu_1_data_master_readdata),                                      //                                                     .readdata
		.cpu_1_data_master_readdatavalid                            (cpu_1_data_master_readdatavalid),                                 //                                                     .readdatavalid
		.cpu_1_data_master_write                                    (cpu_1_data_master_write),                                         //                                                     .write
		.cpu_1_data_master_writedata                                (cpu_1_data_master_writedata),                                     //                                                     .writedata
		.cpu_1_data_master_debugaccess                              (cpu_1_data_master_debugaccess),                                   //                                                     .debugaccess
		.cpu_1_instruction_master_address                           (cpu_1_instruction_master_address),                                //                             cpu_1_instruction_master.address
		.cpu_1_instruction_master_waitrequest                       (cpu_1_instruction_master_waitrequest),                            //                                                     .waitrequest
		.cpu_1_instruction_master_read                              (cpu_1_instruction_master_read),                                   //                                                     .read
		.cpu_1_instruction_master_readdata                          (cpu_1_instruction_master_readdata),                               //                                                     .readdata
		.cpu_1_instruction_master_readdatavalid                     (cpu_1_instruction_master_readdatavalid),                          //                                                     .readdatavalid
		.cpu_0_debug_mem_slave_address                              (mm_interconnect_0_cpu_0_debug_mem_slave_address),                 //                                cpu_0_debug_mem_slave.address
		.cpu_0_debug_mem_slave_write                                (mm_interconnect_0_cpu_0_debug_mem_slave_write),                   //                                                     .write
		.cpu_0_debug_mem_slave_read                                 (mm_interconnect_0_cpu_0_debug_mem_slave_read),                    //                                                     .read
		.cpu_0_debug_mem_slave_readdata                             (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),                //                                                     .readdata
		.cpu_0_debug_mem_slave_writedata                            (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),               //                                                     .writedata
		.cpu_0_debug_mem_slave_byteenable                           (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),              //                                                     .byteenable
		.cpu_0_debug_mem_slave_waitrequest                          (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest),             //                                                     .waitrequest
		.cpu_0_debug_mem_slave_debugaccess                          (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess),             //                                                     .debugaccess
		.cpu_1_debug_mem_slave_address                              (mm_interconnect_0_cpu_1_debug_mem_slave_address),                 //                                cpu_1_debug_mem_slave.address
		.cpu_1_debug_mem_slave_write                                (mm_interconnect_0_cpu_1_debug_mem_slave_write),                   //                                                     .write
		.cpu_1_debug_mem_slave_read                                 (mm_interconnect_0_cpu_1_debug_mem_slave_read),                    //                                                     .read
		.cpu_1_debug_mem_slave_readdata                             (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),                //                                                     .readdata
		.cpu_1_debug_mem_slave_writedata                            (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),               //                                                     .writedata
		.cpu_1_debug_mem_slave_byteenable                           (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),              //                                                     .byteenable
		.cpu_1_debug_mem_slave_waitrequest                          (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest),             //                                                     .waitrequest
		.cpu_1_debug_mem_slave_debugaccess                          (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess),             //                                                     .debugaccess
		.interrupt_counter_0_avalon_slave_0_address                 (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_address),    //                   interrupt_counter_0_avalon_slave_0.address
		.interrupt_counter_0_avalon_slave_0_write                   (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_write),      //                                                     .write
		.interrupt_counter_0_avalon_slave_0_read                    (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_read),       //                                                     .read
		.interrupt_counter_0_avalon_slave_0_readdata                (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_readdata),   //                                                     .readdata
		.interrupt_counter_0_avalon_slave_0_writedata               (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_writedata),  //                                                     .writedata
		.interrupt_counter_0_avalon_slave_0_chipselect              (mm_interconnect_0_interrupt_counter_0_avalon_slave_0_chipselect), //                                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),         //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),           //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),            //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),        //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),       //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),     //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),      //                                                     .chipselect
		.jtag_uart_1_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),         //                        jtag_uart_1_avalon_jtag_slave.address
		.jtag_uart_1_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),           //                                                     .write
		.jtag_uart_1_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),            //                                                     .read
		.jtag_uart_1_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),        //                                                     .readdata
		.jtag_uart_1_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),       //                                                     .writedata
		.jtag_uart_1_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest),     //                                                     .waitrequest
		.jtag_uart_1_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),      //                                                     .chipselect
		.leds_0_s1_address                                          (mm_interconnect_0_leds_0_s1_address),                             //                                            leds_0_s1.address
		.leds_0_s1_write                                            (mm_interconnect_0_leds_0_s1_write),                               //                                                     .write
		.leds_0_s1_readdata                                         (mm_interconnect_0_leds_0_s1_readdata),                            //                                                     .readdata
		.leds_0_s1_writedata                                        (mm_interconnect_0_leds_0_s1_writedata),                           //                                                     .writedata
		.leds_0_s1_chipselect                                       (mm_interconnect_0_leds_0_s1_chipselect),                          //                                                     .chipselect
		.mailbox_simple_0_avmm_msg_receiver_address                 (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address),    //                   mailbox_simple_0_avmm_msg_receiver.address
		.mailbox_simple_0_avmm_msg_receiver_write                   (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write),      //                                                     .write
		.mailbox_simple_0_avmm_msg_receiver_read                    (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read),       //                                                     .read
		.mailbox_simple_0_avmm_msg_receiver_readdata                (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata),   //                                                     .readdata
		.mailbox_simple_0_avmm_msg_receiver_writedata               (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata),  //                                                     .writedata
		.mailbox_simple_0_avmm_msg_sender_address                   (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address),      //                     mailbox_simple_0_avmm_msg_sender.address
		.mailbox_simple_0_avmm_msg_sender_write                     (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write),        //                                                     .write
		.mailbox_simple_0_avmm_msg_sender_read                      (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read),         //                                                     .read
		.mailbox_simple_0_avmm_msg_sender_readdata                  (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata),     //                                                     .readdata
		.mailbox_simple_0_avmm_msg_sender_writedata                 (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata),    //                                                     .writedata
		.mailbox_simple_0_avmm_msg_sender_waitrequest               (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest),  //                                                     .waitrequest
		.mutex_0_s1_address                                         (mm_interconnect_0_mutex_0_s1_address),                            //                                           mutex_0_s1.address
		.mutex_0_s1_write                                           (mm_interconnect_0_mutex_0_s1_write),                              //                                                     .write
		.mutex_0_s1_read                                            (mm_interconnect_0_mutex_0_s1_read),                               //                                                     .read
		.mutex_0_s1_readdata                                        (mm_interconnect_0_mutex_0_s1_readdata),                           //                                                     .readdata
		.mutex_0_s1_writedata                                       (mm_interconnect_0_mutex_0_s1_writedata),                          //                                                     .writedata
		.mutex_0_s1_chipselect                                      (mm_interconnect_0_mutex_0_s1_chipselect),                         //                                                     .chipselect
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                   //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                     //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                  //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),                 //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                     //                                                     .clken
		.onchip_memory2_1_s1_address                                (mm_interconnect_0_onchip_memory2_1_s1_address),                   //                                  onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                                  (mm_interconnect_0_onchip_memory2_1_s1_write),                     //                                                     .write
		.onchip_memory2_1_s1_readdata                               (mm_interconnect_0_onchip_memory2_1_s1_readdata),                  //                                                     .readdata
		.onchip_memory2_1_s1_writedata                              (mm_interconnect_0_onchip_memory2_1_s1_writedata),                 //                                                     .writedata
		.onchip_memory2_1_s1_byteenable                             (mm_interconnect_0_onchip_memory2_1_s1_byteenable),                //                                                     .byteenable
		.onchip_memory2_1_s1_chipselect                             (mm_interconnect_0_onchip_memory2_1_s1_chipselect),                //                                                     .chipselect
		.onchip_memory2_1_s1_clken                                  (mm_interconnect_0_onchip_memory2_1_s1_clken),                     //                                                     .clken
		.perf_count_0_control_slave_address                         (mm_interconnect_0_perf_count_0_control_slave_address),            //                           perf_count_0_control_slave.address
		.perf_count_0_control_slave_write                           (mm_interconnect_0_perf_count_0_control_slave_write),              //                                                     .write
		.perf_count_0_control_slave_readdata                        (mm_interconnect_0_perf_count_0_control_slave_readdata),           //                                                     .readdata
		.perf_count_0_control_slave_writedata                       (mm_interconnect_0_perf_count_0_control_slave_writedata),          //                                                     .writedata
		.perf_count_0_control_slave_begintransfer                   (mm_interconnect_0_perf_count_0_control_slave_begintransfer),      //                                                     .begintransfer
		.perf_count_1_control_slave_address                         (mm_interconnect_0_perf_count_1_control_slave_address),            //                           perf_count_1_control_slave.address
		.perf_count_1_control_slave_write                           (mm_interconnect_0_perf_count_1_control_slave_write),              //                                                     .write
		.perf_count_1_control_slave_readdata                        (mm_interconnect_0_perf_count_1_control_slave_readdata),           //                                                     .readdata
		.perf_count_1_control_slave_writedata                       (mm_interconnect_0_perf_count_1_control_slave_writedata),          //                                                     .writedata
		.perf_count_1_control_slave_begintransfer                   (mm_interconnect_0_perf_count_1_control_slave_begintransfer),      //                                                     .begintransfer
		.timer_0_s1_address                                         (mm_interconnect_0_timer_0_s1_address),                            //                                           timer_0_s1.address
		.timer_0_s1_write                                           (mm_interconnect_0_timer_0_s1_write),                              //                                                     .write
		.timer_0_s1_readdata                                        (mm_interconnect_0_timer_0_s1_readdata),                           //                                                     .readdata
		.timer_0_s1_writedata                                       (mm_interconnect_0_timer_0_s1_writedata),                          //                                                     .writedata
		.timer_0_s1_chipselect                                      (mm_interconnect_0_timer_0_s1_chipselect),                         //                                                     .chipselect
		.timer_1_s1_address                                         (mm_interconnect_0_timer_1_s1_address),                            //                                           timer_1_s1.address
		.timer_1_s1_write                                           (mm_interconnect_0_timer_1_s1_write),                              //                                                     .write
		.timer_1_s1_readdata                                        (mm_interconnect_0_timer_1_s1_readdata),                           //                                                     .readdata
		.timer_1_s1_writedata                                       (mm_interconnect_0_timer_1_s1_writedata),                          //                                                     .writedata
		.timer_1_s1_chipselect                                      (mm_interconnect_0_timer_1_s1_chipselect)                          //                                                     .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_0_irq_irq)                   //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_1_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_0_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_1_debug_reset_request_reset),        // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_1_debug_reset_request_reset),    // reset_in1.reset
		.reset_in2      (cpu_0_debug_reset_request_reset),    // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
