-- soc_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                                 : in    std_logic                     := '0';             --                              clk.clk
		nios_buttons_external_connection_export : in    std_logic_vector(2 downto 0)  := (others => '0'); -- nios_buttons_external_connection.export
		nios_leds_external_connection_export    : out   std_logic_vector(9 downto 0);                     --    nios_leds_external_connection.export
		parallel_port_0_conduit_end_export      : inout std_logic_vector(31 downto 0) := (others => '0'); --      parallel_port_0_conduit_end.export
		pll_0_sdram_clk_clk                     : out   std_logic;                                        --                  pll_0_sdram_clk.clk
		reset_reset_n                           : in    std_logic                     := '0';             --                            reset.reset_n
		sdram_controller_0_wire_addr            : out   std_logic_vector(12 downto 0);                    --          sdram_controller_0_wire.addr
		sdram_controller_0_wire_ba              : out   std_logic_vector(1 downto 0);                     --                                 .ba
		sdram_controller_0_wire_cas_n           : out   std_logic;                                        --                                 .cas_n
		sdram_controller_0_wire_cke             : out   std_logic;                                        --                                 .cke
		sdram_controller_0_wire_cs_n            : out   std_logic;                                        --                                 .cs_n
		sdram_controller_0_wire_dq              : inout std_logic_vector(15 downto 0) := (others => '0'); --                                 .dq
		sdram_controller_0_wire_dqm             : out   std_logic_vector(1 downto 0);                     --                                 .dqm
		sdram_controller_0_wire_ras_n           : out   std_logic;                                        --                                 .ras_n
		sdram_controller_0_wire_we_n            : out   std_logic                                         --                                 .we_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component counter is
		port (
			Clk        : in  std_logic                     := 'X';             -- clk
			Address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			ChipSelect : in  std_logic                     := 'X';             -- chipselect
			Read       : in  std_logic                     := 'X';             -- read
			Write      : in  std_logic                     := 'X';             -- write
			ReadData   : out std_logic_vector(31 downto 0);                    -- readdata
			WriteData  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nReset     : in  std_logic                     := 'X';             -- reset_n
			IRQ        : out std_logic                                         -- irq
		);
	end component counter;

	component soc_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_jtag_uart_0;

	component soc_system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_nios2_gen2_0;

	component soc_system_nios_buttons is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component soc_system_nios_buttons;

	component soc_system_nios_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component soc_system_nios_leds;

	component parallel_port is
		generic (
			N : integer := 32
		);
		port (
			Clk        : in    std_logic                     := 'X';             -- clk
			Address    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			ChipSelect : in    std_logic                     := 'X';             -- chipselect
			Write      : in    std_logic                     := 'X';             -- write
			WriteData  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Read       : in    std_logic                     := 'X';             -- read
			ReadData   : out   std_logic_vector(31 downto 0);                    -- readdata
			nReset     : in    std_logic                     := 'X';             -- reset_n
			ParPort    : inout std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component parallel_port;

	component soc_system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_pll_0;

	component soc_system_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component soc_system_sdram_controller_0;

	component soc_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid;

	component soc_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                             : in  std_logic                     := 'X';             -- clk
			pll_0_outclk0_clk                                         : in  std_logic                     := 'X';             -- clk
			pll_0_outclk1_clk                                         : in  std_logic                     := 'X';             -- clk
			interupt_counter_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                          : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                      : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                             : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                         : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid                    : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                            : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                      : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                   : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest               : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                      : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid             : out std_logic;                                        -- readdatavalid
			interupt_counter_0_avalon_slave_0_address                 : out std_logic_vector(2 downto 0);                     -- address
			interupt_counter_0_avalon_slave_0_write                   : out std_logic;                                        -- write
			interupt_counter_0_avalon_slave_0_read                    : out std_logic;                                        -- read
			interupt_counter_0_avalon_slave_0_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			interupt_counter_0_avalon_slave_0_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			interupt_counter_0_avalon_slave_0_chipselect              : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                  : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                      : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                        : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                         : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                  : out std_logic;                                        -- debugaccess
			nios_buttons_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			nios_buttons_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_leds_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			nios_leds_s1_write                                        : out std_logic;                                        -- write
			nios_leds_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_leds_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			nios_leds_s1_chipselect                                   : out std_logic;                                        -- chipselect
			parallel_port_0_avalon_slave_0_address                    : out std_logic_vector(2 downto 0);                     -- address
			parallel_port_0_avalon_slave_0_write                      : out std_logic;                                        -- write
			parallel_port_0_avalon_slave_0_read                       : out std_logic;                                        -- read
			parallel_port_0_avalon_slave_0_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			parallel_port_0_avalon_slave_0_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			parallel_port_0_avalon_slave_0_chipselect                 : out std_logic;                                        -- chipselect
			sdram_controller_0_s1_address                             : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_0_s1_write                               : out std_logic;                                        -- write
			sdram_controller_0_s1_read                                : out std_logic;                                        -- read
			sdram_controller_0_s1_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_0_s1_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_0_s1_byteenable                          : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_0_s1_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_0_s1_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_0_s1_chipselect                          : out std_logic;                                        -- chipselect
			sysid_control_slave_address                               : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	component soc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_002;

	signal pll_0_outclk0_clk                                               : std_logic;                     -- pll_0:outclk_0 -> [irq_synchronizer_001:receiver_clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, rst_controller_001:clk, sysid:clock]
	signal pll_0_outclk1_clk                                               : std_logic;                     -- pll_0:outclk_1 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, mm_interconnect_0:pll_0_outclk1_clk, nios2_gen2_0:clk, rst_controller_002:clk, sdram_controller_0:clk]
	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(27 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(27 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_interupt_counter_0_avalon_slave_0_chipselect  : std_logic;                     -- mm_interconnect_0:interupt_counter_0_avalon_slave_0_chipselect -> interupt_counter_0:ChipSelect
	signal mm_interconnect_0_interupt_counter_0_avalon_slave_0_readdata    : std_logic_vector(31 downto 0); -- interupt_counter_0:ReadData -> mm_interconnect_0:interupt_counter_0_avalon_slave_0_readdata
	signal mm_interconnect_0_interupt_counter_0_avalon_slave_0_address     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:interupt_counter_0_avalon_slave_0_address -> interupt_counter_0:Address
	signal mm_interconnect_0_interupt_counter_0_avalon_slave_0_read        : std_logic;                     -- mm_interconnect_0:interupt_counter_0_avalon_slave_0_read -> interupt_counter_0:Read
	signal mm_interconnect_0_interupt_counter_0_avalon_slave_0_write       : std_logic;                     -- mm_interconnect_0:interupt_counter_0_avalon_slave_0_write -> interupt_counter_0:Write
	signal mm_interconnect_0_interupt_counter_0_avalon_slave_0_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:interupt_counter_0_avalon_slave_0_writedata -> interupt_counter_0:WriteData
	signal mm_interconnect_0_parallel_port_0_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:parallel_port_0_avalon_slave_0_chipselect -> parallel_port_0:ChipSelect
	signal mm_interconnect_0_parallel_port_0_avalon_slave_0_readdata       : std_logic_vector(31 downto 0); -- parallel_port_0:ReadData -> mm_interconnect_0:parallel_port_0_avalon_slave_0_readdata
	signal mm_interconnect_0_parallel_port_0_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:parallel_port_0_avalon_slave_0_address -> parallel_port_0:Address
	signal mm_interconnect_0_parallel_port_0_avalon_slave_0_read           : std_logic;                     -- mm_interconnect_0:parallel_port_0_avalon_slave_0_read -> parallel_port_0:Read
	signal mm_interconnect_0_parallel_port_0_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:parallel_port_0_avalon_slave_0_write -> parallel_port_0:Write
	signal mm_interconnect_0_parallel_port_0_avalon_slave_0_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:parallel_port_0_avalon_slave_0_writedata -> parallel_port_0:WriteData
	signal mm_interconnect_0_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_nios_leds_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:nios_leds_s1_chipselect -> nios_leds:chipselect
	signal mm_interconnect_0_nios_leds_s1_readdata                         : std_logic_vector(31 downto 0); -- nios_leds:readdata -> mm_interconnect_0:nios_leds_s1_readdata
	signal mm_interconnect_0_nios_leds_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_leds_s1_address -> nios_leds:address
	signal mm_interconnect_0_nios_leds_s1_write                            : std_logic;                     -- mm_interconnect_0:nios_leds_s1_write -> mm_interconnect_0_nios_leds_s1_write:in
	signal mm_interconnect_0_nios_leds_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_leds_s1_writedata -> nios_leds:writedata
	signal mm_interconnect_0_sdram_controller_0_s1_chipselect              : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	signal mm_interconnect_0_sdram_controller_0_s1_readdata                : std_logic_vector(15 downto 0); -- sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	signal mm_interconnect_0_sdram_controller_0_s1_waitrequest             : std_logic;                     -- sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_0_s1_address                 : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	signal mm_interconnect_0_sdram_controller_0_s1_read                    : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_read -> mm_interconnect_0_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_0_s1_byteenable -> mm_interconnect_0_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_0_s1_readdatavalid           : std_logic;                     -- sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_0_s1_write                   : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_write -> mm_interconnect_0_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_sdram_controller_0_s1_writedata               : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	signal mm_interconnect_0_nios_buttons_s1_readdata                      : std_logic_vector(31 downto 0); -- nios_buttons:readdata -> mm_interconnect_0:nios_buttons_s1_readdata
	signal mm_interconnect_0_nios_buttons_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nios_buttons_s1_address -> nios_buttons:address
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                   : std_logic_vector(0 downto 0);  -- interupt_counter_0:IRQ -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                               : std_logic_vector(0 downto 0);  -- jtag_uart_0:av_irq -> irq_synchronizer_001:receiver_irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:interupt_counter_0_reset_sink_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [irq_synchronizer_001:receiver_reset, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_002_reset_out_reset_req                          : std_logic;                     -- rst_controller_002:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_nios_leds_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_nios_leds_s1_write:inv -> nios_leds:write_n
	signal mm_interconnect_0_sdram_controller_0_s1_read_ports_inv          : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_read:inv -> sdram_controller_0:az_rd_n
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv    : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_0_s1_byteenable:inv -> sdram_controller_0:az_be_n
	signal mm_interconnect_0_sdram_controller_0_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_write:inv -> sdram_controller_0:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [interupt_counter_0:nReset, nios_buttons:reset_n, nios_leds:reset_n, parallel_port_0:nReset]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtag_uart_0:rst_n, sysid:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [nios2_gen2_0:reset_n, sdram_controller_0:reset_n]

begin

	interupt_counter_0 : component counter
		port map (
			Clk        => clk_clk,                                                        --            clock.clk
			Address    => mm_interconnect_0_interupt_counter_0_avalon_slave_0_address,    --   avalon_slave_0.address
			ChipSelect => mm_interconnect_0_interupt_counter_0_avalon_slave_0_chipselect, --                 .chipselect
			Read       => mm_interconnect_0_interupt_counter_0_avalon_slave_0_read,       --                 .read
			Write      => mm_interconnect_0_interupt_counter_0_avalon_slave_0_write,      --                 .write
			ReadData   => mm_interconnect_0_interupt_counter_0_avalon_slave_0_readdata,   --                 .readdata
			WriteData  => mm_interconnect_0_interupt_counter_0_avalon_slave_0_writedata,  --                 .writedata
			nReset     => rst_controller_reset_out_reset_ports_inv,                       --       reset_sink.reset_n
			IRQ        => irq_synchronizer_receiver_irq(0)                                -- interrupt_sender.irq
		);

	jtag_uart_0 : component soc_system_jtag_uart_0
		port map (
			clk            => pll_0_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_001_receiver_irq(0)                             --               irq.irq
		);

	nios2_gen2_0 : component soc_system_nios2_gen2_0
		port map (
			clk                                 => pll_0_outclk1_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	nios_buttons : component soc_system_nios_buttons
		port map (
			clk      => clk_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => mm_interconnect_0_nios_buttons_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_nios_buttons_s1_readdata, --                    .readdata
			in_port  => nios_buttons_external_connection_export     -- external_connection.export
		);

	nios_leds : component soc_system_nios_leds
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_nios_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nios_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nios_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nios_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nios_leds_s1_readdata,        --                    .readdata
			out_port   => nios_leds_external_connection_export            -- external_connection.export
		);

	parallel_port_0 : component parallel_port
		generic map (
			N => 32
		)
		port map (
			Clk        => clk_clk,                                                     --          clock.clk
			Address    => mm_interconnect_0_parallel_port_0_avalon_slave_0_address,    -- avalon_slave_0.address
			ChipSelect => mm_interconnect_0_parallel_port_0_avalon_slave_0_chipselect, --               .chipselect
			Write      => mm_interconnect_0_parallel_port_0_avalon_slave_0_write,      --               .write
			WriteData  => mm_interconnect_0_parallel_port_0_avalon_slave_0_writedata,  --               .writedata
			Read       => mm_interconnect_0_parallel_port_0_avalon_slave_0_read,       --               .read
			ReadData   => mm_interconnect_0_parallel_port_0_avalon_slave_0_readdata,   --               .readdata
			nReset     => rst_controller_reset_out_reset_ports_inv,                    --     reset_sink.reset_n
			ParPort    => parallel_port_0_conduit_end_export                           --    conduit_end.export
		);

	pll_0 : component soc_system_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			outclk_1 => pll_0_outclk1_clk,       -- outclk1.clk
			outclk_2 => pll_0_sdram_clk_clk,     -- outclk2.clk
			locked   => open                     -- (terminated)
		);

	sdram_controller_0 : component soc_system_sdram_controller_0
		port map (
			clk            => pll_0_outclk1_clk,                                            --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,                 -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_0_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_0_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_0_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_0_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_0_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_0_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_0_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_0_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_0_wire_we_n                                  --      .export
		);

	sysid : component soc_system_sysid
		port map (
			clock    => pll_0_outclk0_clk,                                --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                             => clk_clk,                                                        --                                           clk_0_clk.clk
			pll_0_outclk0_clk                                         => pll_0_outclk0_clk,                                              --                                       pll_0_outclk0.clk
			pll_0_outclk1_clk                                         => pll_0_outclk1_clk,                                              --                                       pll_0_outclk1.clk
			interupt_counter_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                 -- interupt_counter_0_reset_sink_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset             => rst_controller_001_reset_out_reset,                             --             jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset            => rst_controller_002_reset_out_reset,                             --            nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                          => nios2_gen2_0_data_master_address,                               --                            nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                      => nios2_gen2_0_data_master_waitrequest,                           --                                                    .waitrequest
			nios2_gen2_0_data_master_byteenable                       => nios2_gen2_0_data_master_byteenable,                            --                                                    .byteenable
			nios2_gen2_0_data_master_read                             => nios2_gen2_0_data_master_read,                                  --                                                    .read
			nios2_gen2_0_data_master_readdata                         => nios2_gen2_0_data_master_readdata,                              --                                                    .readdata
			nios2_gen2_0_data_master_readdatavalid                    => nios2_gen2_0_data_master_readdatavalid,                         --                                                    .readdatavalid
			nios2_gen2_0_data_master_write                            => nios2_gen2_0_data_master_write,                                 --                                                    .write
			nios2_gen2_0_data_master_writedata                        => nios2_gen2_0_data_master_writedata,                             --                                                    .writedata
			nios2_gen2_0_data_master_debugaccess                      => nios2_gen2_0_data_master_debugaccess,                           --                                                    .debugaccess
			nios2_gen2_0_instruction_master_address                   => nios2_gen2_0_instruction_master_address,                        --                     nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest               => nios2_gen2_0_instruction_master_waitrequest,                    --                                                    .waitrequest
			nios2_gen2_0_instruction_master_read                      => nios2_gen2_0_instruction_master_read,                           --                                                    .read
			nios2_gen2_0_instruction_master_readdata                  => nios2_gen2_0_instruction_master_readdata,                       --                                                    .readdata
			nios2_gen2_0_instruction_master_readdatavalid             => nios2_gen2_0_instruction_master_readdatavalid,                  --                                                    .readdatavalid
			interupt_counter_0_avalon_slave_0_address                 => mm_interconnect_0_interupt_counter_0_avalon_slave_0_address,    --                   interupt_counter_0_avalon_slave_0.address
			interupt_counter_0_avalon_slave_0_write                   => mm_interconnect_0_interupt_counter_0_avalon_slave_0_write,      --                                                    .write
			interupt_counter_0_avalon_slave_0_read                    => mm_interconnect_0_interupt_counter_0_avalon_slave_0_read,       --                                                    .read
			interupt_counter_0_avalon_slave_0_readdata                => mm_interconnect_0_interupt_counter_0_avalon_slave_0_readdata,   --                                                    .readdata
			interupt_counter_0_avalon_slave_0_writedata               => mm_interconnect_0_interupt_counter_0_avalon_slave_0_writedata,  --                                                    .writedata
			interupt_counter_0_avalon_slave_0_chipselect              => mm_interconnect_0_interupt_counter_0_avalon_slave_0_chipselect, --                                                    .chipselect
			jtag_uart_0_avalon_jtag_slave_address                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,        --                       jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,          --                                                    .write
			jtag_uart_0_avalon_jtag_slave_read                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,           --                                                    .read
			jtag_uart_0_avalon_jtag_slave_readdata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,       --                                                    .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,      --                                                    .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,    --                                                    .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,     --                                                    .chipselect
			nios2_gen2_0_debug_mem_slave_address                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,         --                        nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,           --                                                    .write
			nios2_gen2_0_debug_mem_slave_read                         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,            --                                                    .read
			nios2_gen2_0_debug_mem_slave_readdata                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,        --                                                    .readdata
			nios2_gen2_0_debug_mem_slave_writedata                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,       --                                                    .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,      --                                                    .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,     --                                                    .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,     --                                                    .debugaccess
			nios_buttons_s1_address                                   => mm_interconnect_0_nios_buttons_s1_address,                      --                                     nios_buttons_s1.address
			nios_buttons_s1_readdata                                  => mm_interconnect_0_nios_buttons_s1_readdata,                     --                                                    .readdata
			nios_leds_s1_address                                      => mm_interconnect_0_nios_leds_s1_address,                         --                                        nios_leds_s1.address
			nios_leds_s1_write                                        => mm_interconnect_0_nios_leds_s1_write,                           --                                                    .write
			nios_leds_s1_readdata                                     => mm_interconnect_0_nios_leds_s1_readdata,                        --                                                    .readdata
			nios_leds_s1_writedata                                    => mm_interconnect_0_nios_leds_s1_writedata,                       --                                                    .writedata
			nios_leds_s1_chipselect                                   => mm_interconnect_0_nios_leds_s1_chipselect,                      --                                                    .chipselect
			parallel_port_0_avalon_slave_0_address                    => mm_interconnect_0_parallel_port_0_avalon_slave_0_address,       --                      parallel_port_0_avalon_slave_0.address
			parallel_port_0_avalon_slave_0_write                      => mm_interconnect_0_parallel_port_0_avalon_slave_0_write,         --                                                    .write
			parallel_port_0_avalon_slave_0_read                       => mm_interconnect_0_parallel_port_0_avalon_slave_0_read,          --                                                    .read
			parallel_port_0_avalon_slave_0_readdata                   => mm_interconnect_0_parallel_port_0_avalon_slave_0_readdata,      --                                                    .readdata
			parallel_port_0_avalon_slave_0_writedata                  => mm_interconnect_0_parallel_port_0_avalon_slave_0_writedata,     --                                                    .writedata
			parallel_port_0_avalon_slave_0_chipselect                 => mm_interconnect_0_parallel_port_0_avalon_slave_0_chipselect,    --                                                    .chipselect
			sdram_controller_0_s1_address                             => mm_interconnect_0_sdram_controller_0_s1_address,                --                               sdram_controller_0_s1.address
			sdram_controller_0_s1_write                               => mm_interconnect_0_sdram_controller_0_s1_write,                  --                                                    .write
			sdram_controller_0_s1_read                                => mm_interconnect_0_sdram_controller_0_s1_read,                   --                                                    .read
			sdram_controller_0_s1_readdata                            => mm_interconnect_0_sdram_controller_0_s1_readdata,               --                                                    .readdata
			sdram_controller_0_s1_writedata                           => mm_interconnect_0_sdram_controller_0_s1_writedata,              --                                                    .writedata
			sdram_controller_0_s1_byteenable                          => mm_interconnect_0_sdram_controller_0_s1_byteenable,             --                                                    .byteenable
			sdram_controller_0_s1_readdatavalid                       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,          --                                                    .readdatavalid
			sdram_controller_0_s1_waitrequest                         => mm_interconnect_0_sdram_controller_0_s1_waitrequest,            --                                                    .waitrequest
			sdram_controller_0_s1_chipselect                          => mm_interconnect_0_sdram_controller_0_s1_chipselect,             --                                                    .chipselect
			sysid_control_slave_address                               => mm_interconnect_0_sysid_control_slave_address,                  --                                 sysid_control_slave.address
			sysid_control_slave_readdata                              => mm_interconnect_0_sysid_control_slave_readdata                  --                                                    .readdata
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => pll_0_outclk1_clk,                  --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,                  --       receiver_clk.clk
			sender_clk     => pll_0_outclk1_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                      --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_0_outclk1_clk,                      --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_nios_leds_s1_write_ports_inv <= not mm_interconnect_0_nios_leds_s1_write;

	mm_interconnect_0_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_read;

	mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of soc_system
