-- soc_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                           : in  std_logic                    := '0'; --                        clk.clk
		leds_0_external_connection_export : out std_logic_vector(7 downto 0);        -- leds_0_external_connection.export
		reset_reset_n                     : in  std_logic                    := '0'  --                      reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component soc_system_cpu_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_cpu_0;

	component soc_system_cpu_1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_cpu_1;

	component counter is
		port (
			Clk        : in  std_logic                     := 'X';             -- clk
			IRQ        : out std_logic;                                        -- irq
			nReset     : in  std_logic                     := 'X';             -- reset_n
			Address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			ChipSelect : in  std_logic                     := 'X';             -- chipselect
			Read       : in  std_logic                     := 'X';             -- read
			Write      : in  std_logic                     := 'X';             -- write
			ReadData   : out std_logic_vector(31 downto 0);                    -- readdata
			WriteData  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component counter;

	component soc_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_jtag_uart_0;

	component soc_system_leds_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component soc_system_leds_0;

	component altera_avalon_mailbox is
		generic (
			DWIDTH : integer := 32;
			AWIDTH : integer := 2
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			rst_n                : in  std_logic                     := 'X';             -- reset_n
			avmm_snd_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_snd_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_snd_write       : in  std_logic                     := 'X';             -- write
			avmm_snd_read        : in  std_logic                     := 'X';             -- read
			avmm_snd_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_snd_waitrequest : out std_logic;                                        -- waitrequest
			irq_msg              : out std_logic;                                        -- irq
			avmm_rcv_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read        : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write       : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq_space            : out std_logic                                         -- irq
		);
	end component altera_avalon_mailbox;

	component soc_system_mutex_0 is
		port (
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk           : in  std_logic                     := 'X';             -- clk
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			address       : in  std_logic                     := 'X'              -- address
		);
	end component soc_system_mutex_0;

	component soc_system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component soc_system_onchip_memory2_0;

	component soc_system_onchip_memory2_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component soc_system_onchip_memory2_1;

	component soc_system_perf_count_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component soc_system_perf_count_0;

	component soc_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_timer_0;

	component soc_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			cpu_0_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			cpu_1_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			interrupt_counter_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_0_data_master_address                                  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_0_data_master_waitrequest                              : out std_logic;                                        -- waitrequest
			cpu_0_data_master_byteenable                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_0_data_master_read                                     : in  std_logic                     := 'X';             -- read
			cpu_0_data_master_readdata                                 : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_data_master_readdatavalid                            : out std_logic;                                        -- readdatavalid
			cpu_0_data_master_write                                    : in  std_logic                     := 'X';             -- write
			cpu_0_data_master_writedata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_0_data_master_debugaccess                              : in  std_logic                     := 'X';             -- debugaccess
			cpu_0_instruction_master_address                           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_0_instruction_master_waitrequest                       : out std_logic;                                        -- waitrequest
			cpu_0_instruction_master_read                              : in  std_logic                     := 'X';             -- read
			cpu_0_instruction_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_instruction_master_readdatavalid                     : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_address                                  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_1_data_master_waitrequest                              : out std_logic;                                        -- waitrequest
			cpu_1_data_master_byteenable                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_1_data_master_read                                     : in  std_logic                     := 'X';             -- read
			cpu_1_data_master_readdata                                 : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_data_master_readdatavalid                            : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_write                                    : in  std_logic                     := 'X';             -- write
			cpu_1_data_master_writedata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_1_data_master_debugaccess                              : in  std_logic                     := 'X';             -- debugaccess
			cpu_1_instruction_master_address                           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_1_instruction_master_waitrequest                       : out std_logic;                                        -- waitrequest
			cpu_1_instruction_master_read                              : in  std_logic                     := 'X';             -- read
			cpu_1_instruction_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_instruction_master_readdatavalid                     : out std_logic;                                        -- readdatavalid
			cpu_0_debug_mem_slave_address                              : out std_logic_vector(8 downto 0);                     -- address
			cpu_0_debug_mem_slave_write                                : out std_logic;                                        -- write
			cpu_0_debug_mem_slave_read                                 : out std_logic;                                        -- read
			cpu_0_debug_mem_slave_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_0_debug_mem_slave_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_0_debug_mem_slave_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_0_debug_mem_slave_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			cpu_0_debug_mem_slave_debugaccess                          : out std_logic;                                        -- debugaccess
			cpu_1_debug_mem_slave_address                              : out std_logic_vector(8 downto 0);                     -- address
			cpu_1_debug_mem_slave_write                                : out std_logic;                                        -- write
			cpu_1_debug_mem_slave_read                                 : out std_logic;                                        -- read
			cpu_1_debug_mem_slave_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_1_debug_mem_slave_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_1_debug_mem_slave_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_1_debug_mem_slave_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			cpu_1_debug_mem_slave_debugaccess                          : out std_logic;                                        -- debugaccess
			interrupt_counter_0_avalon_slave_0_address                 : out std_logic_vector(2 downto 0);                     -- address
			interrupt_counter_0_avalon_slave_0_write                   : out std_logic;                                        -- write
			interrupt_counter_0_avalon_slave_0_read                    : out std_logic;                                        -- read
			interrupt_counter_0_avalon_slave_0_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			interrupt_counter_0_avalon_slave_0_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			interrupt_counter_0_avalon_slave_0_chipselect              : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                        : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                         : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   : out std_logic;                                        -- chipselect
			jtag_uart_1_avalon_jtag_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_1_avalon_jtag_slave_write                        : out std_logic;                                        -- write
			jtag_uart_1_avalon_jtag_slave_read                         : out std_logic;                                        -- read
			jtag_uart_1_avalon_jtag_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_1_avalon_jtag_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_1_avalon_jtag_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_1_avalon_jtag_slave_chipselect                   : out std_logic;                                        -- chipselect
			leds_0_s1_address                                          : out std_logic_vector(1 downto 0);                     -- address
			leds_0_s1_write                                            : out std_logic;                                        -- write
			leds_0_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_0_s1_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			leds_0_s1_chipselect                                       : out std_logic;                                        -- chipselect
			mailbox_simple_0_avmm_msg_receiver_address                 : out std_logic_vector(1 downto 0);                     -- address
			mailbox_simple_0_avmm_msg_receiver_write                   : out std_logic;                                        -- write
			mailbox_simple_0_avmm_msg_receiver_read                    : out std_logic;                                        -- read
			mailbox_simple_0_avmm_msg_receiver_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mailbox_simple_0_avmm_msg_receiver_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			mailbox_simple_0_avmm_msg_sender_address                   : out std_logic_vector(1 downto 0);                     -- address
			mailbox_simple_0_avmm_msg_sender_write                     : out std_logic;                                        -- write
			mailbox_simple_0_avmm_msg_sender_read                      : out std_logic;                                        -- read
			mailbox_simple_0_avmm_msg_sender_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mailbox_simple_0_avmm_msg_sender_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			mailbox_simple_0_avmm_msg_sender_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			mutex_0_s1_address                                         : out std_logic_vector(0 downto 0);                     -- address
			mutex_0_s1_write                                           : out std_logic;                                        -- write
			mutex_0_s1_read                                            : out std_logic;                                        -- read
			mutex_0_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mutex_0_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			mutex_0_s1_chipselect                                      : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_address                                : out std_logic_vector(13 downto 0);                    -- address
			onchip_memory2_0_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                  : out std_logic;                                        -- clken
			onchip_memory2_1_s1_address                                : out std_logic_vector(13 downto 0);                    -- address
			onchip_memory2_1_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_1_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_1_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_1_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_1_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_1_s1_clken                                  : out std_logic;                                        -- clken
			perf_count_0_control_slave_address                         : out std_logic_vector(3 downto 0);                     -- address
			perf_count_0_control_slave_write                           : out std_logic;                                        -- write
			perf_count_0_control_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			perf_count_0_control_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			perf_count_0_control_slave_begintransfer                   : out std_logic;                                        -- begintransfer
			perf_count_1_control_slave_address                         : out std_logic_vector(3 downto 0);                     -- address
			perf_count_1_control_slave_write                           : out std_logic;                                        -- write
			perf_count_1_control_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			perf_count_1_control_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			perf_count_1_control_slave_begintransfer                   : out std_logic;                                        -- begintransfer
			timer_0_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                           : out std_logic;                                        -- write
			timer_0_s1_readdata                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                      : out std_logic;                                        -- chipselect
			timer_1_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                                           : out std_logic;                                        -- write
			timer_1_s1_readdata                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                                      : out std_logic                                         -- chipselect
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_002;

	signal cpu_0_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	signal cpu_0_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	signal cpu_0_data_master_debugaccess                                   : std_logic;                     -- cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	signal cpu_0_data_master_address                                       : std_logic_vector(17 downto 0); -- cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	signal cpu_0_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	signal cpu_0_data_master_read                                          : std_logic;                     -- cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	signal cpu_0_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	signal cpu_0_data_master_write                                         : std_logic;                     -- cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	signal cpu_0_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	signal cpu_1_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	signal cpu_1_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	signal cpu_1_data_master_debugaccess                                   : std_logic;                     -- cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	signal cpu_1_data_master_address                                       : std_logic_vector(17 downto 0); -- cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	signal cpu_1_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	signal cpu_1_data_master_read                                          : std_logic;                     -- cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	signal cpu_1_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	signal cpu_1_data_master_write                                         : std_logic;                     -- cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	signal cpu_1_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	signal cpu_1_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	signal cpu_1_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	signal cpu_1_instruction_master_address                                : std_logic_vector(17 downto 0); -- cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	signal cpu_1_instruction_master_read                                   : std_logic;                     -- cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	signal cpu_1_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	signal cpu_0_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	signal cpu_0_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	signal cpu_0_instruction_master_address                                : std_logic_vector(17 downto 0); -- cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	signal cpu_0_instruction_master_read                                   : std_logic;                     -- cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	signal cpu_0_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_interrupt_counter_0_avalon_slave_0_chipselect : std_logic;                     -- mm_interconnect_0:interrupt_counter_0_avalon_slave_0_chipselect -> interrupt_counter_0:ChipSelect
	signal mm_interconnect_0_interrupt_counter_0_avalon_slave_0_readdata   : std_logic_vector(31 downto 0); -- interrupt_counter_0:ReadData -> mm_interconnect_0:interrupt_counter_0_avalon_slave_0_readdata
	signal mm_interconnect_0_interrupt_counter_0_avalon_slave_0_address    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:interrupt_counter_0_avalon_slave_0_address -> interrupt_counter_0:Address
	signal mm_interconnect_0_interrupt_counter_0_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:interrupt_counter_0_avalon_slave_0_read -> interrupt_counter_0:Read
	signal mm_interconnect_0_interrupt_counter_0_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:interrupt_counter_0_avalon_slave_0_write -> interrupt_counter_0:Write
	signal mm_interconnect_0_interrupt_counter_0_avalon_slave_0_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:interrupt_counter_0_avalon_slave_0_writedata -> interrupt_counter_0:WriteData
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata     : std_logic_vector(31 downto 0); -- mailbox_simple_0:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_readdata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest  : std_logic;                     -- mailbox_simple_0:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_address -> mailbox_simple_0:avmm_snd_address
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read         : std_logic;                     -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_read -> mailbox_simple_0:avmm_snd_read
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write        : std_logic;                     -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_write -> mailbox_simple_0:avmm_snd_write
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_writedata -> mailbox_simple_0:avmm_snd_writedata
	signal mm_interconnect_0_perf_count_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- perf_count_0:readdata -> mm_interconnect_0:perf_count_0_control_slave_readdata
	signal mm_interconnect_0_perf_count_0_control_slave_address            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:perf_count_0_control_slave_address -> perf_count_0:address
	signal mm_interconnect_0_perf_count_0_control_slave_begintransfer      : std_logic;                     -- mm_interconnect_0:perf_count_0_control_slave_begintransfer -> perf_count_0:begintransfer
	signal mm_interconnect_0_perf_count_0_control_slave_write              : std_logic;                     -- mm_interconnect_0:perf_count_0_control_slave_write -> perf_count_0:write
	signal mm_interconnect_0_perf_count_0_control_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:perf_count_0_control_slave_writedata -> perf_count_0:writedata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest             : std_logic;                     -- cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_0_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	signal mm_interconnect_0_cpu_0_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_0_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	signal mm_interconnect_0_cpu_0_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                   : std_logic_vector(13 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_mutex_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:mutex_0_s1_chipselect -> mutex_0:chipselect
	signal mm_interconnect_0_mutex_0_s1_readdata                           : std_logic_vector(31 downto 0); -- mutex_0:data_to_cpu -> mm_interconnect_0:mutex_0_s1_readdata
	signal mm_interconnect_0_mutex_0_s1_address                            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mutex_0_s1_address -> mutex_0:address
	signal mm_interconnect_0_mutex_0_s1_read                               : std_logic;                     -- mm_interconnect_0:mutex_0_s1_read -> mutex_0:read
	signal mm_interconnect_0_mutex_0_s1_write                              : std_logic;                     -- mm_interconnect_0:mutex_0_s1_write -> mutex_0:write
	signal mm_interconnect_0_mutex_0_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:mutex_0_s1_writedata -> mutex_0:data_from_cpu
	signal mm_interconnect_0_leds_0_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:leds_0_s1_chipselect -> leds_0:chipselect
	signal mm_interconnect_0_leds_0_s1_readdata                            : std_logic_vector(31 downto 0); -- leds_0:readdata -> mm_interconnect_0:leds_0_s1_readdata
	signal mm_interconnect_0_leds_0_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_0_s1_address -> leds_0:address
	signal mm_interconnect_0_leds_0_s1_write                               : std_logic;                     -- mm_interconnect_0:leds_0_s1_write -> mm_interconnect_0_leds_0_s1_write:in
	signal mm_interconnect_0_leds_0_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_0_s1_writedata -> leds_0:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata   : std_logic_vector(31 downto 0); -- mailbox_simple_0:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_address -> mailbox_simple_0:avmm_rcv_address
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read       : std_logic;                     -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_read -> mailbox_simple_0:avmm_rcv_read
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write      : std_logic;                     -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_write -> mailbox_simple_0:avmm_rcv_write
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_writedata -> mailbox_simple_0:avmm_rcv_writedata
	signal mm_interconnect_0_perf_count_1_control_slave_readdata           : std_logic_vector(31 downto 0); -- perf_count_1:readdata -> mm_interconnect_0:perf_count_1_control_slave_readdata
	signal mm_interconnect_0_perf_count_1_control_slave_address            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:perf_count_1_control_slave_address -> perf_count_1:address
	signal mm_interconnect_0_perf_count_1_control_slave_begintransfer      : std_logic;                     -- mm_interconnect_0:perf_count_1_control_slave_begintransfer -> perf_count_1:begintransfer
	signal mm_interconnect_0_perf_count_1_control_slave_write              : std_logic;                     -- mm_interconnect_0:perf_count_1_control_slave_write -> perf_count_1:write
	signal mm_interconnect_0_perf_count_1_control_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:perf_count_1_control_slave_writedata -> perf_count_1:writedata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest             : std_logic;                     -- cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_1_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	signal mm_interconnect_0_cpu_1_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	signal mm_interconnect_0_cpu_1_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_1_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	signal mm_interconnect_0_cpu_1_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_1_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	signal mm_interconnect_0_onchip_memory2_1_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	signal mm_interconnect_0_onchip_memory2_1_s1_address                   : std_logic_vector(13 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	signal mm_interconnect_0_onchip_memory2_1_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	signal mm_interconnect_0_onchip_memory2_1_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	signal mm_interconnect_0_onchip_memory2_1_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	signal mm_interconnect_0_onchip_memory2_1_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	signal mm_interconnect_0_timer_1_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- timer_0:irq -> irq_mapper:receiver3_irq
	signal cpu_0_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu_0:irq
	signal irq_mapper_001_receiver2_irq                                    : std_logic;                     -- jtag_uart_1:av_irq -> irq_mapper_001:receiver2_irq
	signal irq_mapper_001_receiver3_irq                                    : std_logic;                     -- timer_1:irq -> irq_mapper_001:receiver3_irq
	signal cpu_1_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> cpu_1:irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- interrupt_counter_0:IRQ -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- mailbox_simple_0:irq_msg -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [cpu_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal cpu_0_debug_reset_request_reset                                 : std_logic;                     -- cpu_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in2]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:cpu_1_reset_reset_bridge_in_reset_reset, onchip_memory2_1:reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                     -- rst_controller_001:reset_req -> [cpu_1:reset_req, onchip_memory2_1:reset_req, rst_translator_001:reset_req_in]
	signal cpu_1_debug_reset_request_reset                                 : std_logic;                     -- cpu_1:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:interrupt_counter_0_reset_sink_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_leds_0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_leds_0_s1_write:inv -> leds_0:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read:inv -> jtag_uart_1:av_read_n
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write:inv -> jtag_uart_1:av_write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu_0:reset_n, jtag_uart_0:rst_n, perf_count_0:reset_n, timer_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [cpu_1:reset_n, jtag_uart_1:rst_n, perf_count_1:reset_n, timer_1:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [interrupt_counter_0:nReset, leds_0:reset_n, mailbox_simple_0:rst_n, mutex_0:reset_n]

begin

	cpu_0 : component soc_system_cpu_0
		port map (
			clk                                 => clk_clk,                                             --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_0_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_0_data_master_read,                              --                          .read
			d_readdata                          => cpu_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_0_data_master_write,                             --                          .write
			d_writedata                         => cpu_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_0_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_1 : component soc_system_cpu_1
		port map (
			clk                                 => clk_clk,                                             --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,        --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,              --                          .reset_req
			d_address                           => cpu_1_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_1_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_1_data_master_read,                              --                          .read
			d_readdata                          => cpu_1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_1_data_master_write,                             --                          .write
			d_writedata                         => cpu_1_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_1_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_1_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_1_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_1_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_1_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	interrupt_counter_0 : component counter
		port map (
			Clk        => clk_clk,                                                         --            clock.clk
			IRQ        => irq_mapper_receiver1_irq,                                        -- interrupt_sender.irq
			nReset     => rst_controller_002_reset_out_reset_ports_inv,                    --       reset_sink.reset_n
			Address    => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_address,    --   avalon_slave_0.address
			ChipSelect => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_chipselect, --                 .chipselect
			Read       => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_read,       --                 .read
			Write      => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_write,      --                 .write
			ReadData   => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_readdata,   --                 .readdata
			WriteData  => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_writedata   --                 .writedata
		);

	jtag_uart_0 : component soc_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                         --               irq.irq
		);

	jtag_uart_1 : component soc_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver2_irq                                     --               irq.irq
		);

	leds_0 : component soc_system_leds_0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_leds_0_s1_address,          --                  s1.address
			write_n    => mm_interconnect_0_leds_0_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_0_leds_0_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_0_leds_0_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_0_leds_0_s1_readdata,         --                    .readdata
			out_port   => leds_0_external_connection_export             -- external_connection.export
		);

	mailbox_simple_0 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => clk_clk,                                                        --                   clk.clk
			rst_n                => rst_controller_002_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_receiver0_irq,                                       -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                            --           (terminated)
		);

	mutex_0 : component soc_system_mutex_0
		port map (
			reset_n       => rst_controller_002_reset_out_reset_ports_inv, -- reset.reset_n
			clk           => clk_clk,                                      --   clk.clk
			chipselect    => mm_interconnect_0_mutex_0_s1_chipselect,      --    s1.chipselect
			data_from_cpu => mm_interconnect_0_mutex_0_s1_writedata,       --      .writedata
			read          => mm_interconnect_0_mutex_0_s1_read,            --      .read
			write         => mm_interconnect_0_mutex_0_s1_write,           --      .write
			data_to_cpu   => mm_interconnect_0_mutex_0_s1_readdata,        --      .readdata
			address       => mm_interconnect_0_mutex_0_s1_address(0)       --      .address
		);

	onchip_memory2_0 : component soc_system_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	onchip_memory2_1 : component soc_system_onchip_memory2_1
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_1_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_1_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_1_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_1_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	perf_count_0 : component soc_system_perf_count_0
		port map (
			clk           => clk_clk,                                                    --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                   --         reset.reset_n
			address       => mm_interconnect_0_perf_count_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_perf_count_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_perf_count_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_perf_count_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_perf_count_0_control_slave_writedata      --              .writedata
		);

	perf_count_1 : component soc_system_perf_count_0
		port map (
			clk           => clk_clk,                                                    --           clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,               --         reset.reset_n
			address       => mm_interconnect_0_perf_count_1_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_perf_count_1_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_perf_count_1_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_perf_count_1_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_perf_count_1_control_slave_writedata      --              .writedata
		);

	timer_0 : component soc_system_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                      --   irq.irq
		);

	timer_1 : component soc_system_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_001_receiver3_irq                  --   irq.irq
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                              => clk_clk,                                                         --                                            clk_0_clk.clk
			cpu_0_reset_reset_bridge_in_reset_reset                    => rst_controller_reset_out_reset,                                  --                    cpu_0_reset_reset_bridge_in_reset.reset
			cpu_1_reset_reset_bridge_in_reset_reset                    => rst_controller_001_reset_out_reset,                              --                    cpu_1_reset_reset_bridge_in_reset.reset
			interrupt_counter_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                              -- interrupt_counter_0_reset_sink_reset_bridge_in_reset.reset
			cpu_0_data_master_address                                  => cpu_0_data_master_address,                                       --                                    cpu_0_data_master.address
			cpu_0_data_master_waitrequest                              => cpu_0_data_master_waitrequest,                                   --                                                     .waitrequest
			cpu_0_data_master_byteenable                               => cpu_0_data_master_byteenable,                                    --                                                     .byteenable
			cpu_0_data_master_read                                     => cpu_0_data_master_read,                                          --                                                     .read
			cpu_0_data_master_readdata                                 => cpu_0_data_master_readdata,                                      --                                                     .readdata
			cpu_0_data_master_readdatavalid                            => cpu_0_data_master_readdatavalid,                                 --                                                     .readdatavalid
			cpu_0_data_master_write                                    => cpu_0_data_master_write,                                         --                                                     .write
			cpu_0_data_master_writedata                                => cpu_0_data_master_writedata,                                     --                                                     .writedata
			cpu_0_data_master_debugaccess                              => cpu_0_data_master_debugaccess,                                   --                                                     .debugaccess
			cpu_0_instruction_master_address                           => cpu_0_instruction_master_address,                                --                             cpu_0_instruction_master.address
			cpu_0_instruction_master_waitrequest                       => cpu_0_instruction_master_waitrequest,                            --                                                     .waitrequest
			cpu_0_instruction_master_read                              => cpu_0_instruction_master_read,                                   --                                                     .read
			cpu_0_instruction_master_readdata                          => cpu_0_instruction_master_readdata,                               --                                                     .readdata
			cpu_0_instruction_master_readdatavalid                     => cpu_0_instruction_master_readdatavalid,                          --                                                     .readdatavalid
			cpu_1_data_master_address                                  => cpu_1_data_master_address,                                       --                                    cpu_1_data_master.address
			cpu_1_data_master_waitrequest                              => cpu_1_data_master_waitrequest,                                   --                                                     .waitrequest
			cpu_1_data_master_byteenable                               => cpu_1_data_master_byteenable,                                    --                                                     .byteenable
			cpu_1_data_master_read                                     => cpu_1_data_master_read,                                          --                                                     .read
			cpu_1_data_master_readdata                                 => cpu_1_data_master_readdata,                                      --                                                     .readdata
			cpu_1_data_master_readdatavalid                            => cpu_1_data_master_readdatavalid,                                 --                                                     .readdatavalid
			cpu_1_data_master_write                                    => cpu_1_data_master_write,                                         --                                                     .write
			cpu_1_data_master_writedata                                => cpu_1_data_master_writedata,                                     --                                                     .writedata
			cpu_1_data_master_debugaccess                              => cpu_1_data_master_debugaccess,                                   --                                                     .debugaccess
			cpu_1_instruction_master_address                           => cpu_1_instruction_master_address,                                --                             cpu_1_instruction_master.address
			cpu_1_instruction_master_waitrequest                       => cpu_1_instruction_master_waitrequest,                            --                                                     .waitrequest
			cpu_1_instruction_master_read                              => cpu_1_instruction_master_read,                                   --                                                     .read
			cpu_1_instruction_master_readdata                          => cpu_1_instruction_master_readdata,                               --                                                     .readdata
			cpu_1_instruction_master_readdatavalid                     => cpu_1_instruction_master_readdatavalid,                          --                                                     .readdatavalid
			cpu_0_debug_mem_slave_address                              => mm_interconnect_0_cpu_0_debug_mem_slave_address,                 --                                cpu_0_debug_mem_slave.address
			cpu_0_debug_mem_slave_write                                => mm_interconnect_0_cpu_0_debug_mem_slave_write,                   --                                                     .write
			cpu_0_debug_mem_slave_read                                 => mm_interconnect_0_cpu_0_debug_mem_slave_read,                    --                                                     .read
			cpu_0_debug_mem_slave_readdata                             => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,                --                                                     .readdata
			cpu_0_debug_mem_slave_writedata                            => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,               --                                                     .writedata
			cpu_0_debug_mem_slave_byteenable                           => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,              --                                                     .byteenable
			cpu_0_debug_mem_slave_waitrequest                          => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest,             --                                                     .waitrequest
			cpu_0_debug_mem_slave_debugaccess                          => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess,             --                                                     .debugaccess
			cpu_1_debug_mem_slave_address                              => mm_interconnect_0_cpu_1_debug_mem_slave_address,                 --                                cpu_1_debug_mem_slave.address
			cpu_1_debug_mem_slave_write                                => mm_interconnect_0_cpu_1_debug_mem_slave_write,                   --                                                     .write
			cpu_1_debug_mem_slave_read                                 => mm_interconnect_0_cpu_1_debug_mem_slave_read,                    --                                                     .read
			cpu_1_debug_mem_slave_readdata                             => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,                --                                                     .readdata
			cpu_1_debug_mem_slave_writedata                            => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,               --                                                     .writedata
			cpu_1_debug_mem_slave_byteenable                           => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,              --                                                     .byteenable
			cpu_1_debug_mem_slave_waitrequest                          => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest,             --                                                     .waitrequest
			cpu_1_debug_mem_slave_debugaccess                          => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess,             --                                                     .debugaccess
			interrupt_counter_0_avalon_slave_0_address                 => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_address,    --                   interrupt_counter_0_avalon_slave_0.address
			interrupt_counter_0_avalon_slave_0_write                   => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_write,      --                                                     .write
			interrupt_counter_0_avalon_slave_0_read                    => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_read,       --                                                     .read
			interrupt_counter_0_avalon_slave_0_readdata                => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_readdata,   --                                                     .readdata
			interrupt_counter_0_avalon_slave_0_writedata               => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_writedata,  --                                                     .writedata
			interrupt_counter_0_avalon_slave_0_chipselect              => mm_interconnect_0_interrupt_counter_0_avalon_slave_0_chipselect, --                                                     .chipselect
			jtag_uart_0_avalon_jtag_slave_address                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,         --                        jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,           --                                                     .write
			jtag_uart_0_avalon_jtag_slave_read                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,            --                                                     .read
			jtag_uart_0_avalon_jtag_slave_readdata                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                                                     .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                                                     .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      --                                                     .chipselect
			jtag_uart_1_avalon_jtag_slave_address                      => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address,         --                        jtag_uart_1_avalon_jtag_slave.address
			jtag_uart_1_avalon_jtag_slave_write                        => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write,           --                                                     .write
			jtag_uart_1_avalon_jtag_slave_read                         => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read,            --                                                     .read
			jtag_uart_1_avalon_jtag_slave_readdata                     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata,        --                                                     .readdata
			jtag_uart_1_avalon_jtag_slave_writedata                    => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata,       --                                                     .writedata
			jtag_uart_1_avalon_jtag_slave_waitrequest                  => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest,     --                                                     .waitrequest
			jtag_uart_1_avalon_jtag_slave_chipselect                   => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect,      --                                                     .chipselect
			leds_0_s1_address                                          => mm_interconnect_0_leds_0_s1_address,                             --                                            leds_0_s1.address
			leds_0_s1_write                                            => mm_interconnect_0_leds_0_s1_write,                               --                                                     .write
			leds_0_s1_readdata                                         => mm_interconnect_0_leds_0_s1_readdata,                            --                                                     .readdata
			leds_0_s1_writedata                                        => mm_interconnect_0_leds_0_s1_writedata,                           --                                                     .writedata
			leds_0_s1_chipselect                                       => mm_interconnect_0_leds_0_s1_chipselect,                          --                                                     .chipselect
			mailbox_simple_0_avmm_msg_receiver_address                 => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address,    --                   mailbox_simple_0_avmm_msg_receiver.address
			mailbox_simple_0_avmm_msg_receiver_write                   => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write,      --                                                     .write
			mailbox_simple_0_avmm_msg_receiver_read                    => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read,       --                                                     .read
			mailbox_simple_0_avmm_msg_receiver_readdata                => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata,   --                                                     .readdata
			mailbox_simple_0_avmm_msg_receiver_writedata               => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata,  --                                                     .writedata
			mailbox_simple_0_avmm_msg_sender_address                   => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address,      --                     mailbox_simple_0_avmm_msg_sender.address
			mailbox_simple_0_avmm_msg_sender_write                     => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write,        --                                                     .write
			mailbox_simple_0_avmm_msg_sender_read                      => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read,         --                                                     .read
			mailbox_simple_0_avmm_msg_sender_readdata                  => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata,     --                                                     .readdata
			mailbox_simple_0_avmm_msg_sender_writedata                 => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata,    --                                                     .writedata
			mailbox_simple_0_avmm_msg_sender_waitrequest               => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest,  --                                                     .waitrequest
			mutex_0_s1_address                                         => mm_interconnect_0_mutex_0_s1_address,                            --                                           mutex_0_s1.address
			mutex_0_s1_write                                           => mm_interconnect_0_mutex_0_s1_write,                              --                                                     .write
			mutex_0_s1_read                                            => mm_interconnect_0_mutex_0_s1_read,                               --                                                     .read
			mutex_0_s1_readdata                                        => mm_interconnect_0_mutex_0_s1_readdata,                           --                                                     .readdata
			mutex_0_s1_writedata                                       => mm_interconnect_0_mutex_0_s1_writedata,                          --                                                     .writedata
			mutex_0_s1_chipselect                                      => mm_interconnect_0_mutex_0_s1_chipselect,                         --                                                     .chipselect
			onchip_memory2_0_s1_address                                => mm_interconnect_0_onchip_memory2_0_s1_address,                   --                                  onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                  => mm_interconnect_0_onchip_memory2_0_s1_write,                     --                                                     .write
			onchip_memory2_0_s1_readdata                               => mm_interconnect_0_onchip_memory2_0_s1_readdata,                  --                                                     .readdata
			onchip_memory2_0_s1_writedata                              => mm_interconnect_0_onchip_memory2_0_s1_writedata,                 --                                                     .writedata
			onchip_memory2_0_s1_byteenable                             => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                --                                                     .byteenable
			onchip_memory2_0_s1_chipselect                             => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                --                                                     .chipselect
			onchip_memory2_0_s1_clken                                  => mm_interconnect_0_onchip_memory2_0_s1_clken,                     --                                                     .clken
			onchip_memory2_1_s1_address                                => mm_interconnect_0_onchip_memory2_1_s1_address,                   --                                  onchip_memory2_1_s1.address
			onchip_memory2_1_s1_write                                  => mm_interconnect_0_onchip_memory2_1_s1_write,                     --                                                     .write
			onchip_memory2_1_s1_readdata                               => mm_interconnect_0_onchip_memory2_1_s1_readdata,                  --                                                     .readdata
			onchip_memory2_1_s1_writedata                              => mm_interconnect_0_onchip_memory2_1_s1_writedata,                 --                                                     .writedata
			onchip_memory2_1_s1_byteenable                             => mm_interconnect_0_onchip_memory2_1_s1_byteenable,                --                                                     .byteenable
			onchip_memory2_1_s1_chipselect                             => mm_interconnect_0_onchip_memory2_1_s1_chipselect,                --                                                     .chipselect
			onchip_memory2_1_s1_clken                                  => mm_interconnect_0_onchip_memory2_1_s1_clken,                     --                                                     .clken
			perf_count_0_control_slave_address                         => mm_interconnect_0_perf_count_0_control_slave_address,            --                           perf_count_0_control_slave.address
			perf_count_0_control_slave_write                           => mm_interconnect_0_perf_count_0_control_slave_write,              --                                                     .write
			perf_count_0_control_slave_readdata                        => mm_interconnect_0_perf_count_0_control_slave_readdata,           --                                                     .readdata
			perf_count_0_control_slave_writedata                       => mm_interconnect_0_perf_count_0_control_slave_writedata,          --                                                     .writedata
			perf_count_0_control_slave_begintransfer                   => mm_interconnect_0_perf_count_0_control_slave_begintransfer,      --                                                     .begintransfer
			perf_count_1_control_slave_address                         => mm_interconnect_0_perf_count_1_control_slave_address,            --                           perf_count_1_control_slave.address
			perf_count_1_control_slave_write                           => mm_interconnect_0_perf_count_1_control_slave_write,              --                                                     .write
			perf_count_1_control_slave_readdata                        => mm_interconnect_0_perf_count_1_control_slave_readdata,           --                                                     .readdata
			perf_count_1_control_slave_writedata                       => mm_interconnect_0_perf_count_1_control_slave_writedata,          --                                                     .writedata
			perf_count_1_control_slave_begintransfer                   => mm_interconnect_0_perf_count_1_control_slave_begintransfer,      --                                                     .begintransfer
			timer_0_s1_address                                         => mm_interconnect_0_timer_0_s1_address,                            --                                           timer_0_s1.address
			timer_0_s1_write                                           => mm_interconnect_0_timer_0_s1_write,                              --                                                     .write
			timer_0_s1_readdata                                        => mm_interconnect_0_timer_0_s1_readdata,                           --                                                     .readdata
			timer_0_s1_writedata                                       => mm_interconnect_0_timer_0_s1_writedata,                          --                                                     .writedata
			timer_0_s1_chipselect                                      => mm_interconnect_0_timer_0_s1_chipselect,                         --                                                     .chipselect
			timer_1_s1_address                                         => mm_interconnect_0_timer_1_s1_address,                            --                                           timer_1_s1.address
			timer_1_s1_write                                           => mm_interconnect_0_timer_1_s1_write,                              --                                                     .write
			timer_1_s1_readdata                                        => mm_interconnect_0_timer_1_s1_readdata,                           --                                                     .readdata
			timer_1_s1_writedata                                       => mm_interconnect_0_timer_1_s1_writedata,                          --                                                     .writedata
			timer_1_s1_chipselect                                      => mm_interconnect_0_timer_1_s1_chipselect                          --                                                     .chipselect
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => cpu_0_irq_irq                   --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_001_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_001_receiver3_irq,       -- receiver3.irq
			sender_irq    => cpu_1_irq_irq                       --    sender.irq
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_0_debug_reset_request_reset,    -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => cpu_1_debug_reset_request_reset,        -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_1_debug_reset_request_reset,    -- reset_in1.reset
			reset_in2      => cpu_0_debug_reset_request_reset,    -- reset_in2.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_leds_0_s1_write_ports_inv <= not mm_interconnect_0_leds_0_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of soc_system
